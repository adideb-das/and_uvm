
interface intf();
    // ------------------- port declaration-------------------------------------
    logic   a;
    logic   b;
    logic out;
    //--------------------------------------------------------------------------
endinterface

